module hello;

  initial begin
    $write("Hello, Verilog World!!\n");
  end

endmodule
